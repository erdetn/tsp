// Erdet Nasufi erdet.nasufi@gmail.com Copyrights 2022 (C) //

module tsp

pub fn version() string {
	return '0.1'
}
