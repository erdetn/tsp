module tsp

pub fn version() string {
	return '0.1'
}
